class spi_tran extends uvm_sequence_item;
  //Please fill in the Data Types and Variables.

  `uvm_object_utils(spi_tran)

  function new(string name = "spi_tran");
    super.new(name);
  endfunction
endclass
